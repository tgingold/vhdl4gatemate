library ieee;
use ieee.std_logic_1164.all;
package cc_components is
  component CC_IBUF
    generic (
      PIN_NAME: string := "UNPLACED";
      V_IO: string := "UNDEFINED";
      PULLUP: std_logic_vector (0 downto 0) := "X";
      PULLDOWN: std_logic_vector (0 downto 0) := "X";
      KEEPER: std_logic_vector (0 downto 0) := "X";
      SCHMITT_TRIGGER: std_logic_vector (0 downto 0) := "X";
      DELAY_IBF: std_logic_vector (3 downto 0) := "XXXX";
      FF_IBF: std_logic_vector (0 downto 0) := "X"
    );
    port (
      I: in std_logic;
      Y: out std_logic
    );
  end component;
  component CC_OBUF
    generic (
      PIN_NAME: string := "UNPLACED";
      V_IO: string := "UNDEFINED";
      DRIVE: string := "UNDEFINED";
      SLEW: string := "UNDEFINED";
      DELAY_OBF: std_logic_vector (3 downto 0) := "XXXX";
      FF_OBF: std_logic_vector (0 downto 0) := "X"
    );
    port (
      A: in std_logic;
      O: out std_logic
    );
  end component;
  component CC_TOBUF
    generic (
      PIN_NAME: string := "UNPLACED";
      V_IO: string := "UNDEFINED";
      DRIVE: string := "UNDEFINED";
      SLEW: string := "UNDEFINED";
      PULLUP: std_logic_vector (0 downto 0) := "X";
      PULLDOWN: std_logic_vector (0 downto 0) := "X";
      KEEPER: std_logic_vector (0 downto 0) := "X";
      DELAY_OBF: std_logic_vector (3 downto 0) := "XXXX";
      FF_OBF: std_logic_vector (0 downto 0) := "X"
    );
    port (
      A: in std_logic;
      T: in std_logic;
      O: out std_logic
    );
  end component;
  component CC_IOBUF
    generic (
      PIN_NAME: string := "UNPLACED";
      V_IO: string := "UNDEFINED";
      DRIVE: string := "UNDEFINED";
      SLEW: string := "UNDEFINED";
      PULLUP: std_logic_vector (0 downto 0) := "X";
      PULLDOWN: std_logic_vector (0 downto 0) := "X";
      KEEPER: std_logic_vector (0 downto 0) := "X";
      SCHMITT_TRIGGER: std_logic_vector (0 downto 0) := "X";
      DELAY_IBF: std_logic_vector (3 downto 0) := "XXXX";
      DELAY_OBF: std_logic_vector (3 downto 0) := "XXXX";
      FF_IBF: std_logic_vector (0 downto 0) := "X";
      FF_OBF: std_logic_vector (0 downto 0) := "X"
    );
    port (
      A: in std_logic;
      T: in std_logic;
      Y: out std_logic;
      IO: inout std_logic
    );
  end component;
  component CC_LVDS_IBUF
    generic (
      PIN_NAME_P: string := "UNPLACED";
      PIN_NAME_N: string := "UNPLACED";
      V_IO: string := "UNDEFINED";
      LVDS_RTERM: std_logic_vector (0 downto 0) := "X";
      DELAY_IBF: std_logic_vector (3 downto 0) := "XXXX";
      FF_IBF: std_logic_vector (0 downto 0) := "X"
    );
    port (
      I_P: in std_logic;
      I_N: in std_logic;
      Y: out std_logic
    );
  end component;
  component CC_LVDS_OBUF
    generic (
      PIN_NAME_P: string := "UNPLACED";
      PIN_NAME_N: string := "UNPLACED";
      V_IO: string := "UNDEFINED";
      LVDS_BOOST: std_logic_vector (0 downto 0) := "X";
      DELAY_OBF: std_logic_vector (3 downto 0) := "XXXX";
      FF_OBF: std_logic_vector (0 downto 0) := "X"
    );
    port (
      A: in std_logic;
      O_P: out std_logic;
      O_N: out std_logic
    );
  end component;
  component CC_LVDS_TOBUF
    generic (
      PIN_NAME_P: string := "UNPLACED";
      PIN_NAME_N: string := "UNPLACED";
      V_IO: string := "UNDEFINED";
      LVDS_BOOST: std_logic_vector (0 downto 0) := "X";
      DELAY_OBF: std_logic_vector (3 downto 0) := "XXXX";
      FF_OBF: std_logic_vector (0 downto 0) := "X"
    );
    port (
      A: in std_logic;
      T: in std_logic;
      O_P: out std_logic;
      O_N: out std_logic
    );
  end component;
  component CC_LVDS_IOBUF
    generic (
      PIN_NAME_P: string := "UNPLACED";
      PIN_NAME_N: string := "UNPLACED";
      V_IO: string := "UNDEFINED";
      LVDS_RTERM: std_logic_vector (0 downto 0) := "X";
      LVDS_BOOST: std_logic_vector (0 downto 0) := "X";
      DELAY_IBF: std_logic_vector (3 downto 0) := "XXXX";
      DELAY_OBF: std_logic_vector (3 downto 0) := "XXXX";
      FF_IBF: std_logic_vector (0 downto 0) := "X";
      FF_OBF: std_logic_vector (0 downto 0) := "X"
    );
    port (
      A: in std_logic;
      T: in std_logic;
      IO_P: inout std_logic;
      IO_N: inout std_logic;
      Y: out std_logic
    );
  end component;
  component CC_IDDR
    generic (
      CLK_INV: std_logic_vector (0 downto 0) := "0"
    );
    port (
      D: in std_logic;
      CLK: in std_logic;
      Q0: out string;
      Q1: out std_logic
    );
  end component;
  component CC_ODDR
    generic (
      CLK_INV: std_logic_vector (0 downto 0) := "0"
    );
    port (
      D0: in std_logic;
      D1: in std_logic;
      CLK: in std_logic;
      DDR: in std_logic;
      Q: out std_logic
    );
  end component;
  component CC_DFF
    generic (
      CLK_INV: std_logic_vector (0 downto 0) := "0";
      EN_INV: std_logic_vector (0 downto 0) := "0";
      SR_INV: std_logic_vector (0 downto 0) := "0";
      SR_VAL: std_logic_vector (0 downto 0) := "0";
      INIT: std_logic_vector (0 downto 0) := "X"
    );
    port (
      D: in std_logic;
      CLK: in std_logic;
      EN: in std_logic;
      SR: in std_logic;
      Q: out string
    );
  end component;
  component CC_DLT
    generic (
      G_INV: std_logic_vector (0 downto 0) := "0";
      SR_INV: std_logic_vector (0 downto 0) := "0";
      SR_VAL: std_logic_vector (0 downto 0) := "0";
      INIT: std_logic_vector (0 downto 0) := "X"
    );
    port (
      D: in std_logic;
      G: in std_logic;
      SR: in std_logic;
      Q: out string
    );
  end component;
  component CC_LUT1
    generic (
      INIT: std_logic_vector (1 downto 0) := "00"
    );
    port (
      O: out std_logic;
      I0: in std_logic
    );
  end component;
  component CC_LUT2
    generic (
      INIT: std_logic_vector (3 downto 0) := "0000"
    );
    port (
      O: out std_logic;
      I0: in std_logic;
      I1: in std_logic
    );
  end component;
  component CC_LUT3
    generic (
      INIT: std_logic_vector (7 downto 0) := "00000000"
    );
    port (
      O: out std_logic;
      I0: in std_logic;
      I1: in std_logic;
      I2: in std_logic
    );
  end component;
  component CC_LUT4
    generic (
      INIT: std_logic_vector (15 downto 0) := "0000000000000000"
    );
    port (
      O: out std_logic;
      I0: in std_logic;
      I1: in std_logic;
      I2: in std_logic;
      I3: in std_logic
    );
  end component;
  component CC_MX2
    port (
      D0: in std_logic;
      D1: in std_logic;
      S0: in std_logic;
      Y: out std_logic
    );
  end component;
  component CC_MX4
    port (
      D0: in std_logic;
      D1: in std_logic;
      D2: in std_logic;
      D3: in std_logic;
      S0: in std_logic;
      S1: in std_logic;
      Y: out std_logic
    );
  end component;
  component CC_MX8
    port (
      D0: in std_logic;
      D1: in std_logic;
      D2: in std_logic;
      D3: in std_logic;
      D4: in std_logic;
      D5: in std_logic;
      D6: in std_logic;
      D7: in std_logic;
      S0: in std_logic;
      S1: in std_logic;
      S2: in std_logic;
      Y: out std_logic
    );
  end component;
  component CC_ADDF
    port (
      A: in std_logic;
      B: in std_logic;
      CI: in std_logic;
      CO: out std_logic;
      S: out std_logic
    );
  end component;
  component CC_MULT
    generic (
      A_WIDTH: integer := 0;
      B_WIDTH: integer := 0;
      P_WIDTH: integer := 0
    );
    port (
      A: in std_logic_vector (A_WIDTH - 1 downto 0);
      B: in std_logic_vector (B_WIDTH - 1 downto 0);
      P: out std_logic_vector (P_WIDTH - 1 downto 0)
    );
  end component;
  component CC_BUFG
    port (
      I: in std_logic;
      O: out std_logic
    );
  end component;
  component CC_BRAM_20K
    generic (
      LOC: string := "UNPLACED";
      A_RD_WIDTH: integer := 0;
      B_RD_WIDTH: integer := 0;
      A_WR_WIDTH: integer := 0;
      B_WR_WIDTH: integer := 0;
      RAM_MODE: string := "SDP";
      A_WR_MODE: string := "NO_CHANGE";
      B_WR_MODE: string := "NO_CHANGE";
      A_CLK_INV: integer := 0;
      B_CLK_INV: integer := 0;
      A_EN_INV: integer := 0;
      B_EN_INV: integer := 0;
      A_WE_INV: integer := 0;
      B_WE_INV: integer := 0;
      A_DO_REG: integer := 0;
      B_DO_REG: integer := 0;
      ECC_EN: integer := 0;
      INIT_00: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_01: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_02: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_03: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_04: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_05: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_06: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_07: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_08: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_09: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_10: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_11: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_12: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_13: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_14: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_15: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_16: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_17: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_18: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_19: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_20: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_21: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_22: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_23: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_24: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_25: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_26: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_27: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_28: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_29: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_30: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_31: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_32: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_33: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_34: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_35: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_36: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_37: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_38: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_39: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
    );
    port (
      A_DO: out std_logic_vector (19 downto 0);
      B_DO: out std_logic_vector (19 downto 0);
      ECC_1B_ERR: out std_logic;
      ECC_2B_ERR: out std_logic;
      A_CLK: in std_logic;
      B_CLK: in std_logic;
      A_EN: in std_logic;
      B_EN: in std_logic;
      A_WE: in std_logic;
      B_WE: in std_logic;
      A_ADDR: in std_logic_vector (15 downto 0);
      B_ADDR: in std_logic_vector (15 downto 0);
      A_DI: in std_logic_vector (19 downto 0);
      B_DI: in std_logic_vector (19 downto 0);
      A_BM: in std_logic_vector (19 downto 0);
      B_BM: in std_logic_vector (19 downto 0)
    );
  end component;
  component CC_BRAM_40K
    generic (
      LOC: string := "UNPLACED";
      CAS: string := "NONE";
      A_RD_WIDTH: integer := 0;
      B_RD_WIDTH: integer := 0;
      A_WR_WIDTH: integer := 0;
      B_WR_WIDTH: integer := 0;
      RAM_MODE: string := "SDP";
      A_WR_MODE: string := "NO_CHANGE";
      B_WR_MODE: string := "NO_CHANGE";
      A_CLK_INV: integer := 0;
      B_CLK_INV: integer := 0;
      A_EN_INV: integer := 0;
      B_EN_INV: integer := 0;
      A_WE_INV: integer := 0;
      B_WE_INV: integer := 0;
      A_DO_REG: integer := 0;
      B_DO_REG: integer := 0;
      A_ECC_EN: integer := 0;
      B_ECC_EN: integer := 0;
      INIT_00: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_01: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_02: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_03: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_04: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_05: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_06: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_07: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_08: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_09: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_10: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_11: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_12: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_13: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_14: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_15: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_16: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_17: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_18: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_19: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_20: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_21: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_22: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_23: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_24: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_25: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_26: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_27: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_28: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_29: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_30: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_31: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_32: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_33: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_34: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_35: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_36: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_37: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_38: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_39: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_40: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_41: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_42: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_43: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_44: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_45: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_46: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_47: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_48: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_49: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_4A: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_4B: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_4C: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_4D: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_4E: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_4F: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_50: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_51: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_52: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_53: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_54: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_55: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_56: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_57: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_58: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_59: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_5A: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_5B: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_5C: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_5D: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_5E: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_5F: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_60: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_61: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_62: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_63: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_64: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_65: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_66: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_67: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_68: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_69: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_6A: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_6B: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_6C: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_6D: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_6E: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_6F: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_70: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_71: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_72: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_73: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_74: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_75: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_76: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_77: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_78: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_79: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_7A: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_7B: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_7C: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_7D: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_7E: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      INIT_7F: std_logic_vector (319 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
    );
    port (
      A_DO: out std_logic_vector (39 downto 0);
      B_DO: out std_logic_vector (39 downto 0);
      A_ECC_1B_ERR: out std_logic;
      B_ECC_1B_ERR: out std_logic;
      A_ECC_2B_ERR: out std_logic;
      B_ECC_2B_ERR: out std_logic;
      A_CO: out string;
      B_CO: out string;
      A_CLK: in std_logic;
      B_CLK: in std_logic;
      A_EN: in std_logic;
      B_EN: in std_logic;
      A_WE: in std_logic;
      B_WE: in std_logic;
      A_ADDR: in std_logic_vector (15 downto 0);
      B_ADDR: in std_logic_vector (15 downto 0);
      A_DI: in std_logic_vector (39 downto 0);
      B_DI: in std_logic_vector (39 downto 0);
      A_BM: in std_logic_vector (39 downto 0);
      B_BM: in std_logic_vector (39 downto 0);
      A_CI: in std_logic;
      B_CI: in std_logic
    );
  end component;
  component CC_FIFO_40K
    generic (
      LOC: string := "UNPLACED";
      DYN_STAT_SELECT: integer := 0;
      ALMOST_FULL_OFFSET: std_logic_vector (14 downto 0) := "000000000000000";
      ALMOST_EMPTY_OFFSET: std_logic_vector (14 downto 0) := "000000000000000";
      A_WIDTH: integer := 0;
      B_WIDTH: integer := 0;
      RAM_MODE: string := "TDP";
      FIFO_MODE: string := "SYNC";
      A_CLK_INV: integer := 0;
      B_CLK_INV: integer := 0;
      A_EN_INV: integer := 0;
      B_EN_INV: integer := 0;
      A_WE_INV: integer := 0;
      B_WE_INV: integer := 0;
      A_DO_REG: integer := 0;
      B_DO_REG: integer := 0;
      A_ECC_EN: integer := 0;
      B_ECC_EN: integer := 0
    );
    port (
      A_ECC_1B_ERR: out std_logic;
      B_ECC_1B_ERR: out std_logic;
      A_ECC_2B_ERR: out std_logic;
      B_ECC_2B_ERR: out std_logic;
      A_DO: out std_logic_vector (39 downto 0);
      B_DO: out std_logic_vector (39 downto 0);
      A_CLK: in std_logic;
      A_EN: in std_logic;
      A_DI: in std_logic_vector (39 downto 0);
      B_DI: in std_logic_vector (39 downto 0);
      A_BM: in std_logic_vector (39 downto 0);
      B_BM: in std_logic_vector (39 downto 0);
      B_CLK: in std_logic;
      B_EN: in std_logic;
      B_WE: in std_logic;
      F_RST_N: in std_logic;
      F_ALMOST_FULL_OFFSET: in std_logic_vector (14 downto 0);
      F_ALMOST_EMPTY_OFFSET: in std_logic_vector (14 downto 0);
      F_FULL: out std_logic;
      F_EMPTY: out std_logic;
      F_ALMOST_FULL: out std_logic;
      F_ALMOST_EMPTY: out std_logic;
      F_RD_ERROR: out std_logic;
      F_WR_ERROR: out std_logic;
      F_RD_PTR: out std_logic_vector (15 downto 0);
      F_WR_PTR: out std_logic_vector (15 downto 0)
    );
  end component;
  component CC_L2T4
    generic (
      INIT_L00: std_logic_vector (3 downto 0) := "0000";
      INIT_L01: std_logic_vector (3 downto 0) := "0000";
      INIT_L10: std_logic_vector (3 downto 0) := "0000"
    );
    port (
      O: out std_logic;
      I0: in std_logic;
      I1: in std_logic;
      I2: in std_logic;
      I3: in std_logic
    );
  end component;
  component CC_L2T5
    generic (
      INIT_L02: std_logic_vector (3 downto 0) := "0000";
      INIT_L03: std_logic_vector (3 downto 0) := "0000";
      INIT_L11: std_logic_vector (3 downto 0) := "0000";
      INIT_L20: std_logic_vector (3 downto 0) := "0000"
    );
    port (
      O: out std_logic;
      I0: in std_logic;
      I1: in std_logic;
      I2: in std_logic;
      I3: in std_logic;
      I4: in std_logic
    );
  end component;
  component CC_PLL
    generic (
      REF_CLK: string := "";
      OUT_CLK: string := "";
      PERF_MD: string := "";
      LOCK_REQ: integer := 1;
      CLK270_DOUB: integer := 0;
      CLK180_DOUB: integer := 0;
      LOW_JITTER: integer := 1;
      CI_FILTER_CONST: integer := 2;
      CP_FILTER_CONST: integer := 4
    );
    port (
      CLK_REF: in std_logic;
      CLK_FEEDBACK: in std_logic;
      USR_CLK_REF: in std_logic;
      USR_LOCKED_STDY_RST: in std_logic;
      USR_PLL_LOCKED_STDY: out std_logic;
      USR_PLL_LOCKED: out std_logic;
      CLK270: out std_logic;
      CLK180: out std_logic;
      CLK90: out std_logic;
      CLK0: out std_logic;
      CLK_REF_OUT: out std_logic
    );
  end component;
  component CC_PLL_ADV
    generic (
      PLL_CFG_A: std_logic_vector (95 downto 0) := "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0000000000000000000000000000000000000000000000000000000000000000";
      PLL_CFG_B: std_logic_vector (95 downto 0) := "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0000000000000000000000000000000000000000000000000000000000000000"
    );
    port (
      CLK_REF: in std_logic;
      CLK_FEEDBACK: in std_logic;
      USR_CLK_REF: in std_logic;
      USR_LOCKED_STDY_RST: in std_logic;
      USR_SEL_A_B: in std_logic;
      USR_PLL_LOCKED_STDY: out std_logic;
      USR_PLL_LOCKED: out std_logic;
      CLK270: out std_logic;
      CLK180: out std_logic;
      CLK90: out std_logic;
      CLK0: out std_logic;
      CLK_REF_OUT: out std_logic
    );
  end component;
  component CC_SERDES
    generic (
      RX_BUF_RESET_TIME: std_logic_vector (4 downto 0) := "11000";
      RX_PCS_RESET_TIME: std_logic_vector (4 downto 0) := "11000";
      RX_RESET_TIMER_PRESC: std_logic_vector (4 downto 0) := "00000";
      RX_RESET_DONE_GATE: std_logic_vector (0 downto 0) := "0";
      RX_CDR_RESET_TIME: std_logic_vector (4 downto 0) := "11000";
      RX_EQA_RESET_TIME: std_logic_vector (4 downto 0) := "11000";
      RX_PMA_RESET_TIME: std_logic_vector (4 downto 0) := "11000";
      RX_WAIT_CDR_LOCK: std_logic_vector (0 downto 0) := "1";
      RX_CALIB_EN: std_logic_vector (0 downto 0) := "0";
      RX_CALIB_OVR: std_logic_vector (0 downto 0) := "0";
      RX_CALIB_VAL: std_logic_vector (3 downto 0) := "0000";
      RX_RTERM_VCMSEL: std_logic_vector (2 downto 0) := "001";
      RX_RTERM_PD: std_logic_vector (0 downto 0) := "0";
      RX_EQA_CKP_LF: std_logic_vector (7 downto 0) := "11000101";
      RX_EQA_CKP_HF: std_logic_vector (7 downto 0) := "11000101";
      RX_EQA_CKP_OFFSET: std_logic_vector (7 downto 0) := "10000000";
      RX_EN_EQA: std_logic_vector (0 downto 0) := "0";
      RX_EQA_LOCK_CFG: std_logic_vector (3 downto 0) := "0000";
      RX_TH_MON1: std_logic_vector (4 downto 0) := "00010";
      RX_EN_EQA_EXT_VALUE: std_logic_vector (3 downto 0) := "0000";
      RX_TH_MON2: std_logic_vector (4 downto 0) := "00010";
      RX_TAPW: std_logic_vector (4 downto 0) := "00010";
      RX_AFE_OFFSET: std_logic_vector (4 downto 0) := "00010";
      RX_EQA_CONFIG: std_logic_vector (15 downto 0) := "0000001110000000";
      RX_AFE_PEAK: std_logic_vector (4 downto 0) := "00001";
      RX_AFE_GAIN: std_logic_vector (3 downto 0) := "0001";
      RX_AFE_VCMSEL: std_logic_vector (2 downto 0) := "001";
      RX_CDR_CKP: std_logic_vector (7 downto 0) := "00011111";
      RX_CDR_CKI: std_logic_vector (7 downto 0) := "00000000";
      RX_CDR_TRANS_TH: std_logic_vector (8 downto 0) := "000000010";
      RX_CDR_LOCK_CFG: std_logic_vector (5 downto 0) := "110100";
      RX_CDR_FREQ_ACC: std_logic_vector (14 downto 0) := "000000000000000";
      RX_CDR_PHASE_ACC: std_logic_vector (15 downto 0) := "0000000000000000";
      RX_CDR_SET_ACC_CONFIG: std_logic_vector (1 downto 0) := "00";
      RX_CDR_FORCE_LOCK: std_logic_vector (0 downto 0) := "0";
      RX_ALIGN_MCOMMA_VALUE: std_logic_vector (9 downto 0) := "1100000101";
      RX_MCOMMA_ALIGN_OVR: std_logic_vector (0 downto 0) := "0";
      RX_MCOMMA_ALIGN: std_logic_vector (0 downto 0) := "0";
      RX_ALIGN_PCOMMA_VALUE: std_logic_vector (9 downto 0) := "0011111010";
      RX_PCOMMA_ALIGN_OVR: std_logic_vector (0 downto 0) := "0";
      RX_PCOMMA_ALIGN: std_logic_vector (0 downto 0) := "0";
      RX_ALIGN_COMMA_WORD: std_logic_vector (1 downto 0) := "00";
      RX_ALIGN_COMMA_ENABLE: std_logic_vector (9 downto 0) := "1111111111";
      RX_SLIDE_MODE: std_logic_vector (1 downto 0) := "00";
      RX_COMMA_DETECT_EN_OVR: std_logic_vector (0 downto 0) := "0";
      RX_COMMA_DETECT_EN: std_logic_vector (0 downto 0) := "0";
      RX_SLIDE: std_logic_vector (1 downto 0) := "00";
      RX_EYE_MEAS_EN: std_logic_vector (0 downto 0) := "0";
      RX_EYE_MEAS_CFG: std_logic_vector (14 downto 0) := "000000000000000";
      RX_MON_PH_OFFSET: std_logic_vector (5 downto 0) := "000000";
      RX_EI_BIAS: std_logic_vector (3 downto 0) := "0000";
      RX_EI_BW_SEL: std_logic_vector (3 downto 0) := "0010";
      RX_EN_EI_DETECTOR_OVR: std_logic_vector (0 downto 0) := "0";
      RX_EN_EI_DETECTOR: std_logic_vector (0 downto 0) := "0";
      RX_DATA_SEL: std_logic_vector (0 downto 0) := "0";
      RX_BUF_BYPASS: std_logic_vector (0 downto 0) := "0";
      RX_CLKCOR_USE: std_logic_vector (0 downto 0) := "0";
      RX_CLKCOR_MIN_LAT: std_logic_vector (5 downto 0) := "000001";
      RX_CLKCOR_MAX_LAT: std_logic_vector (5 downto 0) := "111001";
      RX_CLKCOR_SEQ_1_0: std_logic_vector (9 downto 0) := "1110111110";
      RX_CLKCOR_SEQ_1_1: std_logic_vector (9 downto 0) := "1110111110";
      RX_CLKCOR_SEQ_1_2: std_logic_vector (9 downto 0) := "1110111110";
      RX_CLKCOR_SEQ_1_3: std_logic_vector (9 downto 0) := "1110111110";
      RX_PMA_LOOPBACK: std_logic_vector (0 downto 0) := "0";
      RX_PCS_LOOPBACK: std_logic_vector (0 downto 0) := "0";
      RX_DATAPATH_SEL: std_logic_vector (1 downto 0) := "11";
      RX_PRBS_OVR: std_logic_vector (0 downto 0) := "0";
      RX_PRBS_SEL: std_logic_vector (2 downto 0) := "000";
      RX_LOOPBACK_OVR: std_logic_vector (0 downto 0) := "0";
      RX_PRBS_CNT_RESET: std_logic_vector (0 downto 0) := "0";
      RX_POWER_DOWN_OVR: std_logic_vector (0 downto 0) := "0";
      RX_POWER_DOWN_N: std_logic_vector (0 downto 0) := "0";
      RX_RESET_OVR: std_logic_vector (0 downto 0) := "0";
      RX_RESET: std_logic_vector (0 downto 0) := "0";
      RX_PMA_RESET_OVR: std_logic_vector (0 downto 0) := "0";
      RX_PMA_RESET: std_logic_vector (0 downto 0) := "0";
      RX_EQA_RESET_OVR: std_logic_vector (0 downto 0) := "0";
      RX_EQA_RESET: std_logic_vector (0 downto 0) := "0";
      RX_CDR_RESET_OVR: std_logic_vector (0 downto 0) := "0";
      RX_CDR_RESET: std_logic_vector (0 downto 0) := "0";
      RX_PCS_RESET_OVR: std_logic_vector (0 downto 0) := "0";
      RX_PCS_RESET: std_logic_vector (0 downto 0) := "0";
      RX_BUF_RESET_OVR: std_logic_vector (0 downto 0) := "0";
      RX_BUF_RESET: std_logic_vector (0 downto 0) := "0";
      RX_POLARITY_OVR: std_logic_vector (0 downto 0) := "0";
      RX_POLARITY: std_logic_vector (0 downto 0) := "0";
      RX_8B10B_EN_OVR: std_logic_vector (0 downto 0) := "0";
      RX_8B10B_EN: std_logic_vector (0 downto 0) := "0";
      RX_8B10B_BYPASS: std_logic_vector (7 downto 0) := "00000000";
      RX_BYTE_REALIGN: std_logic_vector (0 downto 0) := "0";
      RX_DBG_EN: std_logic_vector (0 downto 0) := "0";
      RX_DBG_SEL: std_logic_vector (1 downto 0) := "00";
      RX_DBG_MODE: std_logic_vector (0 downto 0) := "0";
      RX_DBG_SRAM_DELAY: std_logic_vector (5 downto 0) := "101000";
      RX_DBG_ADDR: std_logic_vector (9 downto 0) := "0000000000";
      RX_DBG_RE: std_logic_vector (0 downto 0) := "0";
      RX_DBG_WE: std_logic_vector (0 downto 0) := "0";
      RX_DBG_DATA: std_logic_vector (19 downto 0) := "00000000000000000000";
      TX_SEL_PRE: std_logic_vector (4 downto 0) := "00000";
      TX_SEL_POST: std_logic_vector (4 downto 0) := "00000";
      TX_AMP: std_logic_vector (4 downto 0) := "11110";
      TX_BRANCH_EN_PRE: std_logic_vector (4 downto 0) := "00000";
      TX_BRANCH_EN_MAIN: std_logic_vector (5 downto 0) := "111111";
      TX_BRANCH_EN_POST: std_logic_vector (4 downto 0) := "00000";
      TX_TAIL_CASCODE: std_logic_vector (2 downto 0) := "001";
      TX_DC_ENABLE: std_logic_vector (6 downto 0) := "1111110";
      TX_DC_OFFSET: std_logic_vector (4 downto 0) := "00000";
      TX_CM_RAISE: std_logic_vector (4 downto 0) := "00000";
      TX_CM_THRESHOLD_0: std_logic_vector (4 downto 0) := "01110";
      TX_CM_THRESHOLD_1: std_logic_vector (4 downto 0) := "00001";
      TX_SEL_PRE_EI: std_logic_vector (4 downto 0) := "00000";
      TX_SEL_POST_EI: std_logic_vector (4 downto 0) := "00000";
      TX_AMP_EI: std_logic_vector (4 downto 0) := "11110";
      TX_BRANCH_EN_PRE_EI: std_logic_vector (4 downto 0) := "00000";
      TX_BRANCH_EN_MAIN_EI: std_logic_vector (5 downto 0) := "111111";
      TX_BRANCH_EN_POST_EI: std_logic_vector (4 downto 0) := "00000";
      TX_TAIL_CASCODE_EI: std_logic_vector (2 downto 0) := "001";
      TX_DC_ENABLE_EI: std_logic_vector (6 downto 0) := "1111110";
      TX_DC_OFFSET_EI: std_logic_vector (4 downto 0) := "00000";
      TX_CM_RAISE_EI: std_logic_vector (4 downto 0) := "00000";
      TX_CM_THRESHOLD_0_EI: std_logic_vector (4 downto 0) := "01110";
      TX_CM_THRESHOLD_1_EI: std_logic_vector (4 downto 0) := "00001";
      TX_SEL_PRE_RXDET: std_logic_vector (4 downto 0) := "00000";
      TX_SEL_POST_RXDET: std_logic_vector (4 downto 0) := "00000";
      TX_AMP_RXDET: std_logic_vector (4 downto 0) := "11110";
      TX_BRANCH_EN_PRE_RXDET: std_logic_vector (4 downto 0) := "00000";
      TX_BRANCH_EN_MAIN_RXDET: std_logic_vector (5 downto 0) := "111111";
      TX_BRANCH_EN_POST_RXDET: std_logic_vector (4 downto 0) := "00000";
      TX_TAIL_CASCODE_RXDET: std_logic_vector (2 downto 0) := "001";
      TX_DC_ENABLE_RXDET: std_logic_vector (6 downto 0) := "1111110";
      TX_DC_OFFSET_RXDET: std_logic_vector (4 downto 0) := "00000";
      TX_CM_RAISE_RXDET: std_logic_vector (4 downto 0) := "00000";
      TX_CM_THRESHOLD_0_RXDET: std_logic_vector (4 downto 0) := "01110";
      TX_CM_THRESHOLD_1_RXDET: std_logic_vector (4 downto 0) := "00001";
      TX_CALIB_EN: std_logic_vector (0 downto 0) := "0";
      TX_CALIB_OVR: std_logic_vector (0 downto 0) := "0";
      TX_CALIB_VAL: std_logic_vector (3 downto 0) := "0000";
      TX_CM_REG_KI: std_logic_vector (7 downto 0) := "00000001";
      TX_CM_SAR_EN: std_logic_vector (0 downto 0) := "0";
      TX_CM_REG_EN: std_logic_vector (0 downto 0) := "1";
      TX_PMA_RESET_TIME: std_logic_vector (4 downto 0) := "11000";
      TX_PCS_RESET_TIME: std_logic_vector (4 downto 0) := "11000";
      TX_PCS_RESET_OVR: std_logic_vector (0 downto 0) := "0";
      TX_PCS_RESET: std_logic_vector (0 downto 0) := "0";
      TX_PMA_RESET_OVR: std_logic_vector (0 downto 0) := "0";
      TX_PMA_RESET: std_logic_vector (0 downto 0) := "0";
      TX_RESET_OVR: std_logic_vector (0 downto 0) := "0";
      TX_RESET: std_logic_vector (0 downto 0) := "0";
      TX_PMA_LOOPBACK: std_logic_vector (1 downto 0) := "00";
      TX_PCS_LOOPBACK: std_logic_vector (0 downto 0) := "0";
      TX_DATAPATH_SEL: std_logic_vector (1 downto 0) := "11";
      TX_PRBS_OVR: std_logic_vector (0 downto 0) := "0";
      TX_PRBS_SEL: std_logic_vector (2 downto 0) := "000";
      TX_PRBS_FORCE_ERR: std_logic_vector (0 downto 0) := "0";
      TX_LOOPBACK_OVR: std_logic_vector (0 downto 0) := "0";
      TX_POWER_DOWN_OVR: std_logic_vector (0 downto 0) := "0";
      TX_POWER_DOWN_N: std_logic_vector (0 downto 0) := "0";
      TX_ELEC_IDLE_OVR: std_logic_vector (0 downto 0) := "0";
      TX_ELEC_IDLE: std_logic_vector (0 downto 0) := "0";
      TX_DETECT_RX_OVR: std_logic_vector (0 downto 0) := "0";
      TX_DETECT_RX: std_logic_vector (0 downto 0) := "0";
      TX_POLARITY_OVR: std_logic_vector (0 downto 0) := "0";
      TX_POLARITY: std_logic_vector (0 downto 0) := "0";
      TX_8B10B_EN_OVR: std_logic_vector (0 downto 0) := "0";
      TX_8B10B_EN: std_logic_vector (0 downto 0) := "0";
      TX_DATA_OVR: std_logic_vector (0 downto 0) := "0";
      TX_DATA_CNT: std_logic_vector (2 downto 0) := "000";
      TX_DATA_VALID: std_logic_vector (0 downto 0) := "0";
      PLL_EN_ADPLL_CTRL: std_logic_vector (0 downto 0) := "0";
      PLL_CONFIG_SEL: std_logic_vector (0 downto 0) := "0";
      PLL_SET_OP_LOCK: std_logic_vector (0 downto 0) := "0";
      PLL_ENFORCE_LOCK: std_logic_vector (0 downto 0) := "0";
      PLL_DISABLE_LOCK: std_logic_vector (0 downto 0) := "0";
      PLL_LOCK_WINDOW: std_logic_vector (0 downto 0) := "1";
      PLL_FAST_LOCK: std_logic_vector (0 downto 0) := "1";
      PLL_SYNC_BYPASS: std_logic_vector (0 downto 0) := "0";
      PLL_PFD_SELECT: std_logic_vector (0 downto 0) := "0";
      PLL_REF_BYPASS: std_logic_vector (0 downto 0) := "0";
      PLL_REF_SEL: std_logic_vector (0 downto 0) := "0";
      PLL_REF_RTERM: std_logic_vector (0 downto 0) := "1";
      PLL_FCNTRL: std_logic_vector (5 downto 0) := "010111";
      PLL_MAIN_DIVSEL: std_logic_vector (5 downto 0) := "110110";
      PLL_OUT_DIVSEL: std_logic_vector (1 downto 0) := "00";
      PLL_CI: std_logic_vector (4 downto 0) := "11000";
      PLL_CP: std_logic_vector (9 downto 0) := "0000101000";
      PLL_AO: std_logic_vector (3 downto 0) := "0000";
      PLL_SCAP: std_logic_vector (2 downto 0) := "000";
      PLL_FILTER_SHIFT: std_logic_vector (1 downto 0) := "01";
      PLL_SAR_LIMIT: std_logic_vector (2 downto 0) := "010";
      PLL_FT: std_logic_vector (10 downto 0) := "00000000010";
      PLL_OPEN_LOOP: std_logic_vector (0 downto 0) := "0";
      PLL_SCAP_AUTO_CAL: std_logic_vector (0 downto 0) := "1";
      PLL_BISC_MODE: std_logic_vector (2 downto 0) := "001";
      PLL_BISC_TIMER_MAX: std_logic_vector (3 downto 0) := "1111";
      PLL_BISC_OPT_DET_IND: std_logic_vector (0 downto 0) := "0";
      PLL_BISC_PFD_SEL: std_logic_vector (0 downto 0) := "0";
      PLL_BISC_DLY_DIR: std_logic_vector (0 downto 0) := "0";
      PLL_BISC_COR_DLY: std_logic_vector (2 downto 0) := "100";
      PLL_BISC_CAL_SIGN: std_logic_vector (0 downto 0) := "0";
      PLL_BISC_CAL_AUTO: std_logic_vector (0 downto 0) := "1";
      PLL_BISC_CP_MIN: std_logic_vector (4 downto 0) := "00100";
      PLL_BISC_CP_MAX: std_logic_vector (4 downto 0) := "01001";
      PLL_BISC_CP_START: std_logic_vector (4 downto 0) := "00110";
      PLL_BISC_DLY_PFD_MON_REF: std_logic_vector (4 downto 0) := "00000";
      PLL_BISC_DLY_PFD_MON_DIV: std_logic_vector (4 downto 0) := "01000";
      SERDES_ENABLE: std_logic_vector (0 downto 0) := "0";
      SERDES_AUTO_INIT: std_logic_vector (0 downto 0) := "0";
      SERDES_TESTMODE: std_logic_vector (0 downto 0) := "0"
    );
    port (
      TX_DATA_I: in std_logic_vector (63 downto 0);
      TX_RESET_I: in std_logic;
      TX_PCS_RESET_I: in std_logic;
      TX_PMA_RESET_I: in std_logic;
      PLL_RESET_I: in std_logic;
      TX_POWER_DOWN_N_I: in std_logic;
      TX_POLARITY_I: in std_logic;
      TX_PRBS_SEL_I: in std_logic_vector (2 downto 0);
      TX_PRBS_FORCE_ERR_I: in std_logic;
      TX_8B10B_EN_I: in std_logic;
      TX_8B10B_BYPASS_I: in std_logic_vector (7 downto 0);
      TX_CHAR_IS_K_I: in std_logic_vector (7 downto 0);
      TX_CHAR_DISPMODE_I: in std_logic_vector (7 downto 0);
      TX_CHAR_DISPVAL_I: in std_logic_vector (7 downto 0);
      TX_ELEC_IDLE_I: in std_logic;
      TX_DETECT_RX_I: in std_logic;
      LOOPBACK_I: in std_logic_vector (2 downto 0);
      TX_CLK_I: in std_logic;
      RX_CLK_I: in std_logic;
      RX_RESET_I: in std_logic;
      RX_PMA_RESET_I: in std_logic;
      RX_EQA_RESET_I: in std_logic;
      RX_CDR_RESET_I: in std_logic;
      RX_PCS_RESET_I: in std_logic;
      RX_BUF_RESET_I: in std_logic;
      RX_POWER_DOWN_N_I: in std_logic;
      RX_POLARITY_I: in std_logic;
      RX_PRBS_SEL_I: in std_logic_vector (2 downto 0);
      RX_PRBS_CNT_RESET_I: in std_logic;
      RX_8B10B_EN_I: in std_logic;
      RX_8B10B_BYPASS_I: in std_logic_vector (7 downto 0);
      RX_EN_EI_DETECTOR_I: in std_logic;
      RX_COMMA_DETECT_EN_I: in std_logic;
      RX_SLIDE_I: in std_logic;
      RX_MCOMMA_ALIGN_I: in std_logic;
      RX_PCOMMA_ALIGN_I: in std_logic;
      REGFILE_CLK_I: in std_logic;
      REGFILE_WE_I: in std_logic;
      REGFILE_EN_I: in std_logic;
      REGFILE_ADDR_I: in std_logic_vector (7 downto 0);
      REGFILE_DI_I: in std_logic_vector (15 downto 0);
      REGFILE_MASK_I: in std_logic_vector (15 downto 0);
      RX_DATA_O: out std_logic_vector (63 downto 0);
      RX_NOT_IN_TABLE_O: out std_logic_vector (7 downto 0);
      RX_CHAR_IS_COMMA_O: out std_logic_vector (7 downto 0);
      RX_CHAR_IS_K_O: out std_logic_vector (7 downto 0);
      RX_DISP_ERR_O: out std_logic_vector (7 downto 0);
      TX_DETECT_RX_DONE_O: out std_logic;
      TX_DETECT_RX_PRESENT_O: out std_logic;
      TX_BUF_ERR_O: out std_logic;
      TX_RESET_DONE_O: out std_logic;
      RX_PRBS_ERR_O: out std_logic;
      RX_BUF_ERR_O: out std_logic;
      RX_BYTE_IS_ALIGNED_O: out std_logic;
      RX_BYTE_REALIGN_O: out std_logic;
      RX_RESET_DONE_O: out std_logic;
      RX_EI_EN_O: out std_logic;
      RX_CLK_O: out std_logic;
      PLL_CLK_O: out std_logic;
      REGFILE_DO_O: out std_logic_vector (15 downto 0);
      REGFILE_RDY_O: out std_logic
    );
  end component;
  component CC_CFG_CTRL
    port (
      DATA: in std_logic_vector (7 downto 0);
      CLK: in std_logic;
      EN: in std_logic;
      RECFG: in std_logic;
      VALID: in std_logic
    );
  end component;
  component CC_USR_RSTN
    port (
      USR_RSTN: out std_logic
    );
  end component;

end;
